/home/VLSI/new/lef/gsclib045_macro.lef