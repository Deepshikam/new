/home/VLSI/new/lef/gsclib045_tech.lef